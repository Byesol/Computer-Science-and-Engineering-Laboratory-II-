`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/04/11 06:02:44
// Design Name: 
// Module Name: hadd_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module hadd_tb;
reg a,b,clk;
wire s,c;

hadd u_hadd(
.a(a), .b(b), .s(s), .c(c)
);
initial begin
    a=1'b0;
    b=1'b1;       
    clk = 0;
end

always clk = #10 ~clk;
always @(posedge clk)begin
    a <= #20 ~a;
    b <= #30 ~b;
   
 end
endmodule
